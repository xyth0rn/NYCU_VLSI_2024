* HW4_0_op.sp
*----------------------------------------------------------------------
* Assumption
* lib = cic018.l/tt/N_18 & P_18
* 1. temp 27
* 2. L=0.18um
*----------------------------------------------------------------------

.lib 'cic018.l'  tt
.temp 27
.option post

*----------------------------------------------------------------------
* Simulation netlist
*----------------------------------------------------------------------
Vg  g   gnd 0.9
Vd  d   gnd 0.9
Vdd ndd gnd 1.8

MN1 d g gnd gnd N_18 W=250n L=900n M=1
MP1 d g ndd ndd p_18 W=250n L=270n M=2

*----------------------------------------------------------------------
* Stimulus
*----------------------------------------------------------------------
.option captab=1 	* nodal capacitance table
.op
.end




*----------------------------------------------------------------------
* Result
*----------------------------------------------------------------------
* HW4_1_0_op.lis
*
* nodal capacitance table 
* node    =    cap
* d       =   1.2573f
* g       =   2.6345f
*
* element  mn1       mp1     
* model    n_18.1    p_18.1  
* id       10.0246u  -10.1859u