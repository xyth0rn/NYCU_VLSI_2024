* HW2_1_1.sp
*----------------------------------------------------------------------
.lib 'cic018.l'  tt
.temp 27
.option post

*----------------------------------------------------------------------
* Simulation netlist
*----------------------------------------------------------------------
Vd  d   gnd 0.9
Vg  g   gnd 0.9
Vdd ndd gnd 1.8

MN1 d g gnd gnd N_18 W=0.25u L=0.18u
MP1 d g ndd ndd P_18 W=0.25u L=0.18u

*----------------------------------------------------------------------
* Stimulus
*----------------------------------------------------------------------
.op
.end