* HW4_1_1_2_dc.sp
*----------------------------------------------------------------------
* Assumption
* lib = cic018.l/tt/N_18 & P_18
* 1. temp 27
* 2. L=0.18um
*----------------------------------------------------------------------

.lib 'cic018.l'  tt
.temp 27
.option post

*----------------------------------------------------------------------
* Simulation netlist
*----------------------------------------------------------------------
Vg  g   gnd 0.9
Vd  d   gnd 0.9
Vdd ndd gnd 1.8

MN1 d g gnd gnd N_18 W=250n L=900n M=1
MP1 d g ndd ndd p_18 W=250n L=270n M=2

*----------------------------------------------------------------------
* Stimulus
*----------------------------------------------------------------------
.option dccap=1
.dc vg 0 1.8 0.01
.meas dc cg find cap(g) at=0.9

.print Cmn1=par("lx18(mn1)")	* https://www.ptt.cc/bbs/comm_and_RF/M.1284928485.A.86F.html
.print Cmp1=par("lx18(mp1)")	* https://bbs.eetop.cn/thread-408732-1-1.html
.end




*----------------------------------------------------------------------
* Result
*----------------------------------------------------------------------
* HW4_1_1_2_dc.ms0
* cg               temper         alter#            
* 2.634e-15        27.0000        1      

* AvanWaves
* HW4_1_1_2_dc.png